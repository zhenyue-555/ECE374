LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_signed.ALL;
use ieee.numeric_std.all;

ENTITY MUL IS

 GENERIC (x : INTEGER := 32;
   y : INTEGER := 32);
 
 PORT(m : IN STD_LOGIC_VECTOR(x - 1 DOWNTO 0);
      q : IN STD_LOGIC_VECTOR(y - 1 DOWNTO 0);
      p : OUT STD_LOGIC_VECTOR(x + y - 1 DOWNTO 0);
    --mul_sel : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    i : IN STD_LOGIC
 );   
END MUL;

ARCHITECTURE behavior OF MUL IS

BEGIN



 PROCESS(m,q) 
 variable Pos1, Neg1, zero:  std_logic_vector(31 downto 0);
 variable Output, Result, Pos2, Neg2: std_logic_vector(63 downto 0);
 variable temp: std_logic;
 
 BEGIN
 
 Pos1 := m;
 Neg1:= (0-m);
 Output := x"0000000000000000";
 Zero := x"00000000";
 Pos2 := x"00000000" & STD_LOGIC_VECTOR(shift_left(unsigned(m),1));
 Neg2 := x"00000000" & STD_LOGIC_VECTOR(shift_left(unsigned(0-m),1));
 

 
 for i in 0 to 15 loop
 
	 
    if(i = 0) then
	    if(q(i*2+1 downto i*2) = "00")then
		    Result(31 downto 0) := Zero;
			 temp := Result(31);
			 
		 elsif(q(i*2+1 downto i*2) = "01")then
		    Result(31 downto 0) := Pos1;
			 temp := Result(31);
			 
		 elsif(q(i*2+1 downto i*2) = "10")then
		    Result := Neg2;
			 temp := Result(32);
			 
		 else
		    Result(31 downto 0) := Neg1;
			 temp := Result(31);
			 
		 end if;

	
	else
	   if(q(i*2+1 downto i*2-1) = "000")then
         Result(31 downto 0) := Zero;
			temp := Result(31);
			
		elsif(q(i*2+1 downto i*2-1)= "001")then
		   Result(31 downto 0) := Pos1;
			temp := Result(31);
		
		elsif(q(i*2+1 downto i*2-1)= "010")then
		   Result(31 downto 0) := Pos1;
			temp := Result(31);

		elsif(q(i*2+1 downto i*2-1) = "011")then
		   Result:= Pos2;
			temp := Result(32);
			
		elsif(q(i*2+1 downto i*2-1) = "100")then
		   Result:= Neg2;			
			temp := Result(32);
			
		elsif(q(i*2+1 downto i*2-1) = "101")then
		   Result(31 downto 0):= Neg1;					 
			temp := Result(31);
			
		elsif(q(i*2+1 downto i*2-1) = "110")then
		   Result(31 downto 0):= Neg1;				 
			temp := Result(31);
			
		elsif(q(i*2+1 downto i*2-1) = "111")then
		   Result(31 downto 0):= Zero;
			temp := Result(31);
			
	   end if;
		
    end if;
	 
	 if(temp = '1')then
	    Result(63 downto 32) := x"FFFFFFFF";
	 else
	    Result(63 downto 32) := x"00000000";
	 end if;
	 
	 Result := STD_LOGIC_VECTOR(shift_left(unsigned(Result),i));
	 
	 Output := Output + Result;
	 
end loop;

   p <= Output;

  
 
  
 END PROCESS;
 
END behavior;